module decoder (
  input  logic [31:0]  fetched_instr_i,
  output logic [1:0]   a_sel_o,
  output logic [2:0]   b_sel_o,
  output logic [4:0]   alu_op_o,
  output logic [2:0]   csr_op_o,
  output logic         csr_we_o,
  output logic         mem_req_o,
  output logic         mem_we_o,
  output logic [2:0]   mem_size_o,
  output logic         gpr_we_o,
  output logic [1:0]   wb_sel_o,
  output logic         illegal_instr_o,
  output logic         branch_o,
  output logic         jal_o,
  output logic         jalr_o,
  output logic         mret_o
);
  import decoder_pkg::*;

//  Для удобства дальнейшего описания модуля, 
//  рекомендуется сперва создать сигналы opcode, 
//  func3, func7 и присвоить им соответствующие биты входного сигнала инструкции.
wire logic [2:0]  funct3 ;
wire logic [6:0]  funct7;
wire logic [6:0] opcode;

assign funct3 = fetched_instr_i[14:12];
assign funct7 = fetched_instr_i[31:25];
assign opcode = fetched_instr_i[6:0];

always_comb begin
    //Внутри блока always_comb до начала блока case можно указать базовые значения для всех выходных сигналов. 
    //Это не то же самое, что вариант default в блоке case. Здесь вы можете описать состояния, которые будут использованы чаще всего, 
    //и в этом случае, присваивание сигналу будет выполняться только в том месте, где появится инструкция, требующая значение этого сигнала, 
    //отличное от базового. пусть все нули
    illegal_instr_o = 1'b0;     //Сигнал о некорректной инструкции	
    mret_o = 1'b0;              //Сигнал об инструкции возврата из прерывания/исключения mret
    jalr_o = 1'b0;              //Сигнал об инструкции безусловного перехода jalr
    jal_o = 1'b0;               //Сигнал об инструкции безусловного перехода jal	
    branch_o = 1'b0;            //Сигнал об инструкции условного перехода	
    wb_sel_o = 2'b00;            //Управляющий сигнал мультиплексора для выбора данных, записываемых в регистровый файл
    alu_op_o = ALU_ADD;         //Операция АЛУ	
    csr_we_o = 1'b0;            //Разрешение на запись в CSR	
    csr_op_o = 3'd0;            //Операция модуля CSR	
    mem_req_o = 1'b0;           //Запрос на доступ к памяти (часть интерфейса памяти)	
    mem_we_o = 1'b0;            //Сигнал разрешения записи в память, «write enable» (при равенстве нулю происходит чтение)
    gpr_we_o = 1'b0;            //Сигнал разрешения записи в регистровый файл
    a_sel_o = 2'd0;             //Управляющий сигнал мультиплексора для выбора первого операнда АЛУ
    b_sel_o = 3'd0;             //Управляющий сигнал мультиплексора для выбора второго операнда АЛУ	
    mem_size_o = 3'd0;          //Управляющий сигнал для выбора размера слова при чтении-записи в память (часть интерфейса памяти)
//#####################################################################################################################################################################################################
    case (opcode)
//#####################################################################################################################################################################################################
        LOAD_OPCODE, STORE_OPCODE: begin
        //LOAD	00000	Записать в rd данные из памяти по адресу rs1+imm
        //STORE	01000	Записать в память по адресу rs1+imm данные из 
            mem_req_o = 1'b1;                                          // разрешаем доступ к памяти
            gpr_we_o = (opcode == LOAD_OPCODE) ? 1'b1 : 1'b0;          // load : gpr_we_o=1                        // store: gpr_we_o= 0               :::разрешение записи в регистровый файл 
            wb_sel_o = (opcode == LOAD_OPCODE) ? 2'b01 : wb_sel_o;     // load :   wb_sel_o =  01                  // wb_sel_o = 00:default            :::выбор данных, записываемых в регистровый файл  
            mem_we_o = (opcode == STORE_OPCODE) ? 1'b1 : 1'b0;         // load :   mem_we_o =  0                   //store: mem_we_o = 1               :::разрешения записи в память
            b_sel_o = (opcode == STORE_OPCODE) ? 3'b101 : 3'b001;      // load :   b_sel_o =  001                  //store: b_sel_o =  b101            :::выбора второго операнда АЛУ	
            
            case(funct3)
                LDST_B, LDST_H, LDST_W, LDST_BU, LDST_HU: mem_size_o = funct3;    // проверка на соответсвия командам размера 
                default: illegal_instr_o = 1'b1;                                  // иначе ошибка операции 
            endcase
        end 
//#####################################################################################################################################################################################################                                                                                  
//        store:                                            store : STORE	01000	Записать в память по адресу rs1+imm данные из rs2	Mem[rs1 + imm] = rs2
//  mem_req_o = 1;                                          1. Запись в память mem_req_o = 1 => доступ к памяти
//  gpr_we_o= 0;                                            2. gpr_we_o = 0 => Сигнал запрета записи в регистровый файл
//  wb_sel_o = 00:default;                                  3. Ставим  wb_sel_o = 00 значит выбираем данные получениие с алу
//  mem_we_o = 1;                                           4. mem_we_o = 1 => Сигнал разрешения записи в память
//  b_sel_o =  101;                                         5. тип получаемого imm : b_sel_o = 101 => {[31:25],[11:7]}  -s тип на мультиплексоре
//      ::DEFAULT::                                          
//  alu_op_o = ALU_ADD;                                     6. тип операции alu_op_o = ALU_ADD - значит скложение [rs1 + imm]= mem_adr_0
//  a_sel_o = 2'd0;                                         7. получение a a_sel_o = 2'd0 - c rd1 - по адрессу : 19:15 биты команды
//  mem_size_o = 3'd0;                                      8. Ставим размер записываемого mem_size_o = 3'd0 
// получается записываем в память по адрессу [rs1 + imm]                                                                                      
//#####################################################################################################################################################################################################
//    Load:                                                 store : LOAD	00000	Записать в rd данные из памяти по адресу rs1+imm	rd = Mem[rs1 + imm]
//mem_req_o = 1;                                            1. Запись в память mem_req_o = 1 => доступ к памяти
//gpr_we_o= 1;                                              2. gpr_we_o = 1 => Сигнал разрешения записи в регистровый файл
//wb_sel_o = 01;                                            3. Ставим  wb_sel_o = 01 значит выбираем данные получениие считанные из внешней памяти 
//mem_we_o = 0;                                             4. mem_we_o = 0 => Сигнал запрета записи в память
//b_sel_o =  001;                                           5. тип получаемого imm : b_sel_o = 001 => [31:20]  -I тип на мультиплексоре
//  ::DEFAULT::                                          
//alu_op_o = ALU_ADD;                                      6. тип операции alu_op_o = ALU_ADD - значит скложение [rs1 + imm]= mem_adr_0
//a_sel_o = 2'd0;                                          7. получение a a_sel_o = 2'd0 - c rd1 - по адрессу : 19:15 биты команды
//mem_size_o = 3'd0;                                       8. Ставим размер записываемого mem_size_o = 3'd0 
// получается записываем из памяти по адрессу [rs1 + imm]  в rd по адрессу 11:07 биты команды
//#####################################################################################################################################################################################################
        OP_IMM_OPCODE, OP_OPCODE: begin
            gpr_we_o = 1'b1;
            alu_op_o = funct3;
            case(funct3)
                ALU_ADD, ALU_SLTS, ALU_SLTU, ALU_XOR, ALU_OR, ALU_AND: alu_op_o = funct3;
                default: illegal_instr_o = 1'b1;
            endcase
        end
//#####################################################################################################################################################################################################
//                                                          OP	01100	Записать в rd результат вычисления АЛУ над rs1 и rs2
//  gpr_we_o = 1'b1;                                        1.  gpr_we_o = 1 => Сигнал разрешения записи в регистровый файл
//  alu_op_o = funct3;                                      2.  alu_op_o = funct3; => просто выбор операции которая будет на алу
//     ::DEFAULT::
//  wb_sel_o = 2'b00                                        3.  wb_sel_o = 2'b00;    значит выбираем данные получениие с алу
//  mem_req_o = 1'b0;                                       4.  Запись в память mem_req_o = 0 => доступ к памяти - закрыт
//  mem_we_o = 1'b0;                                        5.  mem_we_o = 0 => Сигнал запрета записи в память
//  a_sel_o = 2'd0;                                         6.  a_sel_o = 2'd0 => данные с RD1 - находящегося по адрессу [19:15] из инструкции
//  b_sel_o = 3'd0;                                         7.  b_sel_o = 3'd0 => данные с RD2 - находящегося по адрессу [24:20] из инструкции
      // то есть мы берем данные с первого регистра и второго реистр по адрессу из инструкции делаем операцию переданую по алуоп и записываем в регистрный файл по адрессу [11:7]
//#####################################################################################################################################################################################################
        AUIPC_OPCODE: begin
            a_sel_o = 2'd1;
            b_sel_o = 3'd2;
            gpr_we_o = 1'b1;
        end
//#####################################################################################################################################################################################################
//                                                          AUIPC	00101	Записать в rd результат сложения непосредственного операнда U-типа imm_u и счетчика команд
//  a_sel_o = 2'd1;                                         1.  a_sel_o = 2'd1 => данные со счетчика команд 
//  b_sel_o = 3'd2;                                         2.  b_sel_o = 3'd2 => тип получаемого imm  => {[31:12],12'h000}  -U тип на мультиплексоре
//  gpr_we_o = 1'b1;                                        3.  gpr_we_o = 1 => Сигнал разрешения записи в регистровый файл
//     ::DEFAULT::
//  alu_op_o = ALU_ADD;                                     4.  тип операции alu_op_o = ALU_ADD - значит скложение [rs1 + imm]= mem_adr_0
//  wb_sel_o = 2'b00                                        5.  wb_sel_o = 2'b00;    значит выбираем данные получениие с алу
//  mem_req_o = 1'b0;                                       6.  Запись в память mem_req_o = 0 => доступ к памяти - закрыт
//  mem_we_o = 1'b0;                                        7.  mem_we_o = 0 => Сигнал запрета записи в память

      // то есть мы берем данные с счетчика команд и складываем с константой смещенной на 12 т.е адресс страницы и записываем в регистрный файл по адрессу [11:7] из инструкции

//#####################################################################################################################################################################################################
        BRANCH_OPCODE: begin
//        localparam ALU_LTS  = 5'b11100;  // Less Than Signed                      FUNCT3<----100 
//        localparam ALU_LTU  = 5'b11110;  // Less Than Unsigned                    FUNCT3<----110
//        localparam ALU_GES  = 5'b11101;  // Great [or] Equal signed               FUNCT3<----101    
//        localparam ALU_GEU  = 5'b11111;  // Great [or] Equal unsigned             FUNCT3<----111    
//        localparam ALU_EQ   = 5'b11000;  // Equal                                 FUNCT3<----000
//        localparam ALU_NE   = 5'b11001;  // Not Equal                             FUNCT3<----001    
            alu_op_o = {2'b11, funct3};   
            branch_o = 1'b1;  
        end
//#####################################################################################################################################################################################################   
//                                                          BRANCH	11000	Увеличить счетчик команд на значение imm, если верен результат сравнения rs1 и rs2
//  alu_op_o = {2'b11, funct3};                             1. alu_op_o = funct3; => просто выбор операции которая будет на алу  
//  branch_o = 1'b1;                                        2. branch_o = 1'b1 => будем прыгать если да и след команда если нет
//  ::DEFAULT::
//  wb_sel_o = 2'b00;                                       3.  wb_sel_o = 2'b00;    значит выбираем данные получениие с алу                
//  mem_req_o = 1'b0;                                       4.  Запись в память mem_req_o = 0 => доступ к памяти - закрыт
//  mem_we_o = 1'b0;                                        5.  mem_we_o = 0 => Сигнал запрета записи в память
//  gpr_we_o = 1'b0;                                        6.  gpr_we_o = 0 => Сигнал запрета записи в регистровый файл
//  a_sel_o = 2'd0;                                         7.  a_sel_o = 2'd0 => данные с RD1 - находящегося по адрессу [19:15] из инструкции
//  b_sel_o = 3'd0;                                         8.  b_sel_o = 3'd0 => данные с RD2 - находящегося по адрессу [24:20] из инструкции
// тут понятно что прыжок либо происходит и тогда прыгает на собранную по частям imm:
//[31] – старший бит смещения (знак)
//[30:25] – старшие биты
//[11:8] – средние биты
//[7] – младший бит
//[0] – всегда 0 (смещение кратно 2)
//#####################################################################################################################################################################################################   
        JALR_OPCODE: begin
          // 
            a_sel_o = 2'd1;    
            b_sel_o = 3'd4; 
            gpr_we_o = 1'b1; 
            jalr_o = 1'b1; 
        end
//#####################################################################################################################################################################################################   
//                                                          JALR	11001	Записать в rd следующий адрес счетчика команд, в счетчик команд записать rs1+imm
//  a_sel_o = 2'd1;                                         1.  a_sel_o = 2'd1 =>данные со счетчика команд 
//  b_sel_o = 3'd4;                                         2.  b_sel_o = 3'd4 => просто константа 4 
//  gpr_we_o = 1'b1;                                        3.  gpr_we_o= 1'b0  => Сигнал разрешений записи в регистровый файл
//  jalr_o = 1'b0;                                          4.  jalr_o = 1'b0 => Сигнал об инструкции безусловного перехода jalr
//  ::DEFAULT::
//  alu_op_o = ALU_ADD;                                     5. тип операции alu_op_o = ALU_ADD - значит скложение [rs1 + imm]= mem_adr_0
//  branch_o = 1'b0;                                        6. branch_o = 1'b0 => переход не условный
//  wb_sel_o = 2'b00;                                       7.  wb_sel_o = 2'b00;    значит выбираем данные получениие с алу                
//  mem_req_o = 1'b0;                                       8.  Запись в память mem_req_o = 0 => доступ к памяти - закрыт
//  mem_we_o = 1'b0;                                        9.  mem_we_o = 0 => Сигнал запрета записи в память
// тут понятно что прыжок происходит на собранную по частям imm+rd1- находящуюся по адрессу[19:15] битах команды, а в rd = pc + 4 или же по адрессу[11:07] битах команды, т.е. след команда
//#####################################################################################################################################################################################################
        JAL_OPCODE: begin
            a_sel_o = 2'd1;
            b_sel_o = 3'd4; 
            gpr_we_o = 1'b1;
            jal_o = 1'b1;
        end
//#####################################################################################################################################################################################################  
        SYSTEM_OPCODE: begin
            case(funct3)
                3'b000: begin
                    case(fetched_instr_i[31:7])
                        25'b001100000010_00000_000_00000: mret_o = 1'b1;
                        default: illegal_instr_o = 1'b1;
                    endcase
                end
                3'b001, 3'b010, 3'b011, 3'b101, 3'b110, 3'b111: begin
                    csr_op_o = funct3;
                    csr_we_o = 1'b1;
                    gpr_we_o = 1'b1;
                    wb_sel_o = 2'd2;
                end
                default: illegal_instr_o = 1'b1;
            endcase
        end
//#####################################################################################################################################################################################################
        default: illegal_instr_o = 1'b1; //если ничего из опкодов не совпало
    endcase
end

endmodule


