module decoder_mega (
  input  logic [31:0]  fetched_instr_i,
  output logic [1:0]   a_sel_o,
  output logic [2:0]   b_sel_o,
  output logic [4:0]   alu_op_o,
  output logic [2:0]   csr_op_o,
  output logic         csr_we_o,
  output logic         mem_req_o,
  output logic         mem_we_o,
  output logic [2:0]   mem_size_o,
  output logic         gpr_we_o,
  output logic [1:0]   wb_sel_o,
  output logic         illegal_instr_o,
  output logic         branch_o,
  output logic         jal_o,
  output logic         jalr_o,
  output logic         mret_o
);
  import decoder_pkg::*;

//  Для удобства дальнейшего описания модуля, 
//  рекомендуется сперва создать сигналы opcode, 
//  func3, func7 и присвоить им соответствующие биты входного сигнала инструкции.
wire logic [2:0]  funct3 ;
wire logic [6:0]  funct7;
wire logic [6:0] opcode;

assign funct3 = fetched_instr_i[14:12];
assign funct7 = fetched_instr_i[31:25];
assign opcode = fetched_instr_i[6:0];

  always_comb begin
 //Проверка на то что 2 младших бита opcode равны '11'
    if(fetched_instr_i[1:0]) begin
    
     //Определение значение по умолчанию
     //Внутри блока always_comb до начала блока case можно указать базовые значения для всех выходных сигналов. 
    //Это не то же самое, что вариант default в блоке case. Здесь вы можете описать состояния, которые будут использованы чаще всего, 
    //и в этом случае, присваивание сигналу будет выполняться только в том месте, где появится инструкция, требующая значение этого сигнала, 
    //отличное от базового. пусть все нули
    illegal_instr_o = 1'b0;     //Сигнал о некорректной инструкции	
    mret_o = 1'b0;              //Сигнал об инструкции возврата из прерывания/исключения mret
    jalr_o = 1'b0;              //Сигнал об инструкции безусловного перехода jalr
    jal_o = 1'b0;               //Сигнал об инструкции безусловного перехода jal	
    branch_o = 1'b0;            //Сигнал об инструкции условного перехода	
    wb_sel_o = 2'b00;            //Управляющий сигнал мультиплексора для выбора данных, записываемых в регистровый файл
    alu_op_o = ALU_ADD;         //Операция АЛУ	
    csr_we_o = 1'b0;            //Разрешение на запись в CSR	
    csr_op_o = 3'd0;            //Операция модуля CSR	
    mem_req_o = 1'b0;           //Запрос на доступ к памяти (часть интерфейса памяти)	
    mem_we_o = 1'b0;            //Сигнал разрешения записи в память, «write enable» (при равенстве нулю происходит чтение)
    gpr_we_o = 1'b0;            //Сигнал разрешения записи в регистровый файл
    a_sel_o = 2'd0;             //Управляющий сигнал мультиплексора для выбора первого операнда АЛУ
    b_sel_o = 3'd0;             //Управляющий сигнал мультиплексора для выбора второго операнда АЛУ	
    mem_size_o = 3'd0;          //Управляющий сигнал для выбора размера слова при чтении-записи в память (часть интерфейса памяти)
 //#####################################################################################################################################################################################################
    case (opcode)
//#####################################################################################################################################################################################################
STORE_OPCODE: begin
          mem_req_o = 1;
          gpr_we_o = 0;
          mem_we_o = 1;
          b_sel_o = OP_B_IMM_S;
         case(funct3)
                LDST_B, LDST_H, LDST_W: mem_size_o = funct3;    // проверка на соответсвия командам размера 

            default : begin illegal_instr_o = 1;  mem_req_o = 0; mem_we_o = 0; end
          endcase
        end
//#####################################################################################################################################################################################################                                                                                  
//        store:                                            store : STORE	01000	Записать в память по адресу rs1+imm данные из rs2	Mem[rs1 + imm] = rs2
//  mem_req_o = 1;                                          1. Запись в память mem_req_o = 1 => доступ к памяти
//  gpr_we_o= 0;                                            2. gpr_we_o = 0 => Сигнал запрета записи в регистровый файл
//  wb_sel_o = 00:default;                                  3. Ставим  wb_sel_o = 00 значит выбираем данные получениие с алу
//  mem_we_o = 1;                                           4. mem_we_o = 1 => Сигнал разрешения записи в память
//  b_sel_o =  OP_B_IMM_S;                                  5. тип получаемого imm : b_sel_o = OP_B_IMM_S => {[31:25],[11:7]}  -s тип на мультиплексоре
//      ::DEFAULT::                                          
//  alu_op_o = ALU_ADD;                                     6. тип операции alu_op_o = ALU_ADD - значит скложение [rs1 + imm]= mem_adr_0
//  a_sel_o = 2'd0;                                         7. получение a a_sel_o = 2'd0 - c rd1 - по адрессу : 19:15 биты команды
//  mem_size_o = 3'd0;                                      8. Ставим размер записываемого mem_size_o = 3'd0 
// получается записываем в память по адрессу [rs1 + imm]                                                                                      
//#####################################################################################################################################################################################################
 LOAD_OPCODE: begin
          mem_req_o = 1;
          gpr_we_o = 1;
          wb_sel_o = 1;
          b_sel_o = OP_B_IMM_I;
          case(funct3)
                LDST_B, LDST_H, LDST_W, LDST_BU, LDST_HU: mem_size_o = funct3;    // проверка на соответсвия командам размера 
                default: illegal_instr_o = 1'b1; mem_req_o = 0; gpr_we_o = 0;;    // иначе ошибка операции  запрет на изменения
            endcase
        end 
//#####################################################################################################################################################################################################
//    Load:                                                 store : LOAD	00000	Записать в rd данные из памяти по адресу rs1+imm	rd = Mem[rs1 + imm]
//mem_req_o = 1;                                            1. Запись в память mem_req_o = 1 => доступ к памяти
//gpr_we_o= 1;                                              2. gpr_we_o = 1 => Сигнал разрешения записи в регистровый файл
//wb_sel_o = 01;                                            3. Ставим  wb_sel_o = 01 значит выбираем данные получениие считанные из внешней памяти 
//mem_we_o = 0;                                             4. mem_we_o = 0 => Сигнал запрета записи в память
//b_sel_o =  OP_B_IMM_I;                                    5. тип получаемого imm : b_sel_o = OP_B_IMM_I => [31:20]  -I тип на мультиплексоре
//  ::DEFAULT::                                          
//alu_op_o = ALU_ADD;                                       6. тип операции alu_op_o = ALU_ADD - значит скложение [rs1 + imm]= mem_adr_0
//a_sel_o = 2'd0;                                           7. получение a a_sel_o = 2'd0 - c rd1 - по адрессу : 19:15 биты команды
//mem_size_o = 3'd0;                                        8. Ставим размер записываемого mem_size_o = 3'd0 
// получается записываем из памяти по адрессу [rs1 + imm]  в rd по адрессу 11:07 биты команды
//#####################################################################################################################################################################################################

      
    end
    else begin 
      illegal_instr_o = 1; 
    end
end
endmodule



